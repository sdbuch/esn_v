// esn7e_demo.v

// Generated using ACDS version 13.1 162 at 2016.08.02.13:56:40

`timescale 1 ps / 1 ps
module esn7e_demo (
		input  wire       clk_clk,            //         clk.clk
		input  wire       reset_reset_n,      //       reset.reset_n
		input  wire       esn_ext_rst_reset,  // esn_ext_rst.reset
		output wire       clk1_locked_export, // clk1_locked.export
		output wire [7:0] led_g_export        //       led_g.export
	);

	wire         altpll_esn_c0_clk;                                                // altpll_esn:c0 -> [EchoStateNetwork_7Units_Expanded_0:clk, avalon_st_adapter:in_clk_0_clk, esn_output_fifo:wrclock, esn_reset_gate:clk]
	wire         esn_reset_gate_reset_out_reset;                                   // esn_reset_gate:reset_out -> [EchoStateNetwork_7Units_Expanded_0:reset, avalon_st_adapter:in_rst_0_reset, esn_output_fifo:wrreset_n]
	wire         nios2_qsys_instruction_master_waitrequest;                        // mm_interconnect_0:nios2_qsys_instruction_master_waitrequest -> nios2_qsys:i_waitrequest
	wire  [19:0] nios2_qsys_instruction_master_address;                            // nios2_qsys:i_address -> mm_interconnect_0:nios2_qsys_instruction_master_address
	wire         nios2_qsys_instruction_master_read;                               // nios2_qsys:i_read -> mm_interconnect_0:nios2_qsys_instruction_master_read
	wire  [31:0] nios2_qsys_instruction_master_readdata;                           // mm_interconnect_0:nios2_qsys_instruction_master_readdata -> nios2_qsys:i_readdata
	wire         nios2_qsys_instruction_master_readdatavalid;                      // mm_interconnect_0:nios2_qsys_instruction_master_readdatavalid -> nios2_qsys:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;        // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;          // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;            // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;         // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;              // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;               // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;           // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire  [31:0] mm_interconnect_0_altpll_esn_pll_slave_writedata;                 // mm_interconnect_0:altpll_esn_pll_slave_writedata -> altpll_esn:writedata
	wire   [1:0] mm_interconnect_0_altpll_esn_pll_slave_address;                   // mm_interconnect_0:altpll_esn_pll_slave_address -> altpll_esn:address
	wire         mm_interconnect_0_altpll_esn_pll_slave_write;                     // mm_interconnect_0:altpll_esn_pll_slave_write -> altpll_esn:write
	wire         mm_interconnect_0_altpll_esn_pll_slave_read;                      // mm_interconnect_0:altpll_esn_pll_slave_read -> altpll_esn:read
	wire  [31:0] mm_interconnect_0_altpll_esn_pll_slave_readdata;                  // altpll_esn:readdata -> mm_interconnect_0:altpll_esn_pll_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_control_slave_address;               // mm_interconnect_0:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire  [31:0] mm_interconnect_0_sysid_qsys_control_slave_readdata;              // sysid_qsys:readdata -> mm_interconnect_0:sysid_qsys_control_slave_readdata
	wire  [31:0] mm_interconnect_0_esn_output_fifo_out_csr_writedata;              // mm_interconnect_0:esn_output_fifo_out_csr_writedata -> esn_output_fifo:rdclk_control_slave_writedata
	wire   [2:0] mm_interconnect_0_esn_output_fifo_out_csr_address;                // mm_interconnect_0:esn_output_fifo_out_csr_address -> esn_output_fifo:rdclk_control_slave_address
	wire         mm_interconnect_0_esn_output_fifo_out_csr_write;                  // mm_interconnect_0:esn_output_fifo_out_csr_write -> esn_output_fifo:rdclk_control_slave_write
	wire         mm_interconnect_0_esn_output_fifo_out_csr_read;                   // mm_interconnect_0:esn_output_fifo_out_csr_read -> esn_output_fifo:rdclk_control_slave_read
	wire  [31:0] mm_interconnect_0_esn_output_fifo_out_csr_readdata;               // esn_output_fifo:rdclk_control_slave_readdata -> mm_interconnect_0:esn_output_fifo_out_csr_readdata
	wire         mm_interconnect_0_nios2_qsys_jtag_debug_module_waitrequest;       // nios2_qsys:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_qsys_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_nios2_qsys_jtag_debug_module_writedata;         // mm_interconnect_0:nios2_qsys_jtag_debug_module_writedata -> nios2_qsys:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_nios2_qsys_jtag_debug_module_address;           // mm_interconnect_0:nios2_qsys_jtag_debug_module_address -> nios2_qsys:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_qsys_jtag_debug_module_write;             // mm_interconnect_0:nios2_qsys_jtag_debug_module_write -> nios2_qsys:jtag_debug_module_write
	wire         mm_interconnect_0_nios2_qsys_jtag_debug_module_read;              // mm_interconnect_0:nios2_qsys_jtag_debug_module_read -> nios2_qsys:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_nios2_qsys_jtag_debug_module_readdata;          // nios2_qsys:jtag_debug_module_readdata -> mm_interconnect_0:nios2_qsys_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_qsys_jtag_debug_module_debugaccess;       // mm_interconnect_0:nios2_qsys_jtag_debug_module_debugaccess -> nios2_qsys:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_nios2_qsys_jtag_debug_module_byteenable;        // mm_interconnect_0:nios2_qsys_jtag_debug_module_byteenable -> nios2_qsys:jtag_debug_module_byteenable
	wire         mm_interconnect_0_esn_output_fifo_out_waitrequest;                // esn_output_fifo:avalonmm_read_slave_waitrequest -> mm_interconnect_0:esn_output_fifo_out_waitrequest
	wire   [0:0] mm_interconnect_0_esn_output_fifo_out_address;                    // mm_interconnect_0:esn_output_fifo_out_address -> esn_output_fifo:avalonmm_read_slave_address
	wire         mm_interconnect_0_esn_output_fifo_out_read;                       // mm_interconnect_0:esn_output_fifo_out_read -> esn_output_fifo:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_esn_output_fifo_out_readdata;                   // esn_output_fifo:avalonmm_read_slave_readdata -> mm_interconnect_0:esn_output_fifo_out_readdata
	wire  [31:0] mm_interconnect_0_led_g_s1_writedata;                             // mm_interconnect_0:led_g_s1_writedata -> led_g:writedata
	wire   [1:0] mm_interconnect_0_led_g_s1_address;                               // mm_interconnect_0:led_g_s1_address -> led_g:address
	wire         mm_interconnect_0_led_g_s1_chipselect;                            // mm_interconnect_0:led_g_s1_chipselect -> led_g:chipselect
	wire         mm_interconnect_0_led_g_s1_write;                                 // mm_interconnect_0:led_g_s1_write -> led_g:write_n
	wire  [31:0] mm_interconnect_0_led_g_s1_readdata;                              // led_g:readdata -> mm_interconnect_0:led_g_s1_readdata
	wire         nios2_qsys_data_master_waitrequest;                               // mm_interconnect_0:nios2_qsys_data_master_waitrequest -> nios2_qsys:d_waitrequest
	wire  [31:0] nios2_qsys_data_master_writedata;                                 // nios2_qsys:d_writedata -> mm_interconnect_0:nios2_qsys_data_master_writedata
	wire  [19:0] nios2_qsys_data_master_address;                                   // nios2_qsys:d_address -> mm_interconnect_0:nios2_qsys_data_master_address
	wire         nios2_qsys_data_master_write;                                     // nios2_qsys:d_write -> mm_interconnect_0:nios2_qsys_data_master_write
	wire         nios2_qsys_data_master_read;                                      // nios2_qsys:d_read -> mm_interconnect_0:nios2_qsys_data_master_read
	wire  [31:0] nios2_qsys_data_master_readdata;                                  // mm_interconnect_0:nios2_qsys_data_master_readdata -> nios2_qsys:d_readdata
	wire         nios2_qsys_data_master_debugaccess;                               // nios2_qsys:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_data_master_debugaccess
	wire         nios2_qsys_data_master_readdatavalid;                             // mm_interconnect_0:nios2_qsys_data_master_readdatavalid -> nios2_qsys:d_readdatavalid
	wire   [3:0] nios2_qsys_data_master_byteenable;                                // nios2_qsys:d_byteenable -> mm_interconnect_0:nios2_qsys_data_master_byteenable
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_writedata;                    // mm_interconnect_0:onchip_memory2_s1_writedata -> onchip_memory2:writedata
	wire  [15:0] mm_interconnect_0_onchip_memory2_s1_address;                      // mm_interconnect_0:onchip_memory2_s1_address -> onchip_memory2:address
	wire         mm_interconnect_0_onchip_memory2_s1_chipselect;                   // mm_interconnect_0:onchip_memory2_s1_chipselect -> onchip_memory2:chipselect
	wire         mm_interconnect_0_onchip_memory2_s1_clken;                        // mm_interconnect_0:onchip_memory2_s1_clken -> onchip_memory2:clken
	wire         mm_interconnect_0_onchip_memory2_s1_write;                        // mm_interconnect_0:onchip_memory2_s1_write -> onchip_memory2:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_readdata;                     // onchip_memory2:readdata -> mm_interconnect_0:onchip_memory2_s1_readdata
	wire   [3:0] mm_interconnect_0_onchip_memory2_s1_byteenable;                   // mm_interconnect_0:onchip_memory2_s1_byteenable -> onchip_memory2:byteenable
	wire         irq_mapper_receiver0_irq;                                         // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                         // esn_output_fifo:rdclk_control_slave_irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_qsys_d_irq_irq;                                             // irq_mapper:sender_irq -> nios2_qsys:d_irq
	wire         echostatenetwork_7units_expanded_0_avalon_streaming_source_valid; // EchoStateNetwork_7Units_Expanded_0:data_valid -> avalon_st_adapter:in_0_valid
	wire  [31:0] echostatenetwork_7units_expanded_0_avalon_streaming_source_data;  // EchoStateNetwork_7Units_Expanded_0:data_out -> avalon_st_adapter:in_0_data
	wire         avalon_st_adapter_out_0_valid;                                    // avalon_st_adapter:out_0_valid -> esn_output_fifo:avalonst_sink_valid
	wire  [31:0] avalon_st_adapter_out_0_data;                                     // avalon_st_adapter:out_0_data -> esn_output_fifo:avalonst_sink_data
	wire         avalon_st_adapter_out_0_ready;                                    // esn_output_fifo:avalonst_sink_ready -> avalon_st_adapter:out_0_ready
	wire         rst_controller_reset_out_reset;                                   // rst_controller:reset_out -> [altpll_esn:reset, esn_output_fifo:rdreset_n, irq_mapper:reset, jtag_uart:rst_n, led_g:reset_n, mm_interconnect_0:nios2_qsys_reset_n_reset_bridge_in_reset_reset, nios2_qsys:reset_n, onchip_memory2:reset, rst_translator:in_reset, sysid_qsys:reset_n]
	wire         rst_controller_reset_out_reset_req;                               // rst_controller:reset_req -> [nios2_qsys:reset_req, onchip_memory2:reset_req, rst_translator:reset_req_in]
	wire         nios2_qsys_jtag_debug_module_reset_reset;                         // nios2_qsys:jtag_debug_module_resetrequest -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	wire         rst_controller_001_reset_out_reset;                               // rst_controller_001:reset_out -> esn_reset_gate:reset_in0

	esn7e_demo_altpll_esn altpll_esn (
		.clk       (clk_clk),                                          //       inclk_interface.clk
		.reset     (rst_controller_reset_out_reset),                   // inclk_interface_reset.reset
		.read      (mm_interconnect_0_altpll_esn_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_altpll_esn_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_altpll_esn_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_altpll_esn_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_altpll_esn_pll_slave_writedata), //                      .writedata
		.c0        (altpll_esn_c0_clk),                                //                    c0.clk
		.areset    (),                                                 //        areset_conduit.export
		.locked    (clk1_locked_export),                               //        locked_conduit.export
		.phasedone ()                                                  //     phasedone_conduit.export
	);

	esn7e_st_src echostatenetwork_7units_expanded_0 (
		.clk        (altpll_esn_c0_clk),                                                //                   clock.clk
		.reset      (esn_reset_gate_reset_out_reset),                                   //                   reset.reset
		.data_valid (echostatenetwork_7units_expanded_0_avalon_streaming_source_valid), // avalon_streaming_source.valid
		.data_out   (echostatenetwork_7units_expanded_0_avalon_streaming_source_data)   //                        .data
	);

	esn7e_demo_nios2_qsys nios2_qsys (
		.clk                                   (clk_clk),                                                    //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                            //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                             (nios2_qsys_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_qsys_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_qsys_data_master_read),                                //                          .read
		.d_readdata                            (nios2_qsys_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_qsys_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_qsys_data_master_write),                               //                          .write
		.d_writedata                           (nios2_qsys_data_master_writedata),                           //                          .writedata
		.d_readdatavalid                       (nios2_qsys_data_master_readdatavalid),                       //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_qsys_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_qsys_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_qsys_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_qsys_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (nios2_qsys_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (nios2_qsys_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_qsys_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_qsys_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_qsys_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_qsys_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_qsys_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_qsys_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_qsys_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_qsys_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_qsys_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                            // custom_instruction_master.readra
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) esn_reset_gate (
		.reset_in0      (rst_controller_001_reset_out_reset), // reset_in0.reset
		.reset_in1      (esn_ext_rst_reset),                  // reset_in1.reset
		.clk            (altpll_esn_c0_clk),                  //       clk.clk
		.reset_out      (esn_reset_gate_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	esn7e_demo_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	esn7e_demo_onchip_memory2 onchip_memory2 (
		.clk        (clk_clk),                                        //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                 // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)              //       .reset_req
	);

	esn7e_demo_sysid_qsys sysid_qsys (
		.clock    (clk_clk),                                             //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                     //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_control_slave_address)   //              .address
	);

	esn7e_demo_led_g led_g (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_led_g_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_g_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_g_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_g_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_g_s1_readdata),   //                    .readdata
		.out_port   (led_g_export)                           // external_connection.export
	);

	esn7e_demo_esn_output_fifo esn_output_fifo (
		.wrclock                         (altpll_esn_c0_clk),                                   //    clk_in.clk
		.wrreset_n                       (~esn_reset_gate_reset_out_reset),                     //  reset_in.reset_n
		.rdclock                         (clk_clk),                                             //   clk_out.clk
		.rdreset_n                       (~rst_controller_reset_out_reset),                     // reset_out.reset_n
		.avalonst_sink_valid             (avalon_st_adapter_out_0_valid),                       //        in.valid
		.avalonst_sink_data              (avalon_st_adapter_out_0_data),                        //          .data
		.avalonst_sink_ready             (avalon_st_adapter_out_0_ready),                       //          .ready
		.avalonmm_read_slave_readdata    (mm_interconnect_0_esn_output_fifo_out_readdata),      //       out.readdata
		.avalonmm_read_slave_read        (mm_interconnect_0_esn_output_fifo_out_read),          //          .read
		.avalonmm_read_slave_address     (mm_interconnect_0_esn_output_fifo_out_address),       //          .address
		.avalonmm_read_slave_waitrequest (mm_interconnect_0_esn_output_fifo_out_waitrequest),   //          .waitrequest
		.rdclk_control_slave_address     (mm_interconnect_0_esn_output_fifo_out_csr_address),   //   out_csr.address
		.rdclk_control_slave_read        (mm_interconnect_0_esn_output_fifo_out_csr_read),      //          .read
		.rdclk_control_slave_writedata   (mm_interconnect_0_esn_output_fifo_out_csr_writedata), //          .writedata
		.rdclk_control_slave_write       (mm_interconnect_0_esn_output_fifo_out_csr_write),     //          .write
		.rdclk_control_slave_readdata    (mm_interconnect_0_esn_output_fifo_out_csr_readdata),  //          .readdata
		.rdclk_control_slave_irq         (irq_mapper_receiver1_irq)                             //   out_irq.irq
	);

	esn7e_demo_mm_interconnect_0 mm_interconnect_0 (
		.clk_50_clk_clk                                 (clk_clk),                                                    //                               clk_50_clk.clk
		.nios2_qsys_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                             // nios2_qsys_reset_n_reset_bridge_in_reset.reset
		.nios2_qsys_data_master_address                 (nios2_qsys_data_master_address),                             //                   nios2_qsys_data_master.address
		.nios2_qsys_data_master_waitrequest             (nios2_qsys_data_master_waitrequest),                         //                                         .waitrequest
		.nios2_qsys_data_master_byteenable              (nios2_qsys_data_master_byteenable),                          //                                         .byteenable
		.nios2_qsys_data_master_read                    (nios2_qsys_data_master_read),                                //                                         .read
		.nios2_qsys_data_master_readdata                (nios2_qsys_data_master_readdata),                            //                                         .readdata
		.nios2_qsys_data_master_readdatavalid           (nios2_qsys_data_master_readdatavalid),                       //                                         .readdatavalid
		.nios2_qsys_data_master_write                   (nios2_qsys_data_master_write),                               //                                         .write
		.nios2_qsys_data_master_writedata               (nios2_qsys_data_master_writedata),                           //                                         .writedata
		.nios2_qsys_data_master_debugaccess             (nios2_qsys_data_master_debugaccess),                         //                                         .debugaccess
		.nios2_qsys_instruction_master_address          (nios2_qsys_instruction_master_address),                      //            nios2_qsys_instruction_master.address
		.nios2_qsys_instruction_master_waitrequest      (nios2_qsys_instruction_master_waitrequest),                  //                                         .waitrequest
		.nios2_qsys_instruction_master_read             (nios2_qsys_instruction_master_read),                         //                                         .read
		.nios2_qsys_instruction_master_readdata         (nios2_qsys_instruction_master_readdata),                     //                                         .readdata
		.nios2_qsys_instruction_master_readdatavalid    (nios2_qsys_instruction_master_readdatavalid),                //                                         .readdatavalid
		.altpll_esn_pll_slave_address                   (mm_interconnect_0_altpll_esn_pll_slave_address),             //                     altpll_esn_pll_slave.address
		.altpll_esn_pll_slave_write                     (mm_interconnect_0_altpll_esn_pll_slave_write),               //                                         .write
		.altpll_esn_pll_slave_read                      (mm_interconnect_0_altpll_esn_pll_slave_read),                //                                         .read
		.altpll_esn_pll_slave_readdata                  (mm_interconnect_0_altpll_esn_pll_slave_readdata),            //                                         .readdata
		.altpll_esn_pll_slave_writedata                 (mm_interconnect_0_altpll_esn_pll_slave_writedata),           //                                         .writedata
		.esn_output_fifo_out_address                    (mm_interconnect_0_esn_output_fifo_out_address),              //                      esn_output_fifo_out.address
		.esn_output_fifo_out_read                       (mm_interconnect_0_esn_output_fifo_out_read),                 //                                         .read
		.esn_output_fifo_out_readdata                   (mm_interconnect_0_esn_output_fifo_out_readdata),             //                                         .readdata
		.esn_output_fifo_out_waitrequest                (mm_interconnect_0_esn_output_fifo_out_waitrequest),          //                                         .waitrequest
		.esn_output_fifo_out_csr_address                (mm_interconnect_0_esn_output_fifo_out_csr_address),          //                  esn_output_fifo_out_csr.address
		.esn_output_fifo_out_csr_write                  (mm_interconnect_0_esn_output_fifo_out_csr_write),            //                                         .write
		.esn_output_fifo_out_csr_read                   (mm_interconnect_0_esn_output_fifo_out_csr_read),             //                                         .read
		.esn_output_fifo_out_csr_readdata               (mm_interconnect_0_esn_output_fifo_out_csr_readdata),         //                                         .readdata
		.esn_output_fifo_out_csr_writedata              (mm_interconnect_0_esn_output_fifo_out_csr_writedata),        //                                         .writedata
		.jtag_uart_avalon_jtag_slave_address            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),      //              jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),        //                                         .write
		.jtag_uart_avalon_jtag_slave_read               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),         //                                         .read
		.jtag_uart_avalon_jtag_slave_readdata           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),     //                                         .readdata
		.jtag_uart_avalon_jtag_slave_writedata          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),    //                                         .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),  //                                         .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),   //                                         .chipselect
		.led_g_s1_address                               (mm_interconnect_0_led_g_s1_address),                         //                                 led_g_s1.address
		.led_g_s1_write                                 (mm_interconnect_0_led_g_s1_write),                           //                                         .write
		.led_g_s1_readdata                              (mm_interconnect_0_led_g_s1_readdata),                        //                                         .readdata
		.led_g_s1_writedata                             (mm_interconnect_0_led_g_s1_writedata),                       //                                         .writedata
		.led_g_s1_chipselect                            (mm_interconnect_0_led_g_s1_chipselect),                      //                                         .chipselect
		.nios2_qsys_jtag_debug_module_address           (mm_interconnect_0_nios2_qsys_jtag_debug_module_address),     //             nios2_qsys_jtag_debug_module.address
		.nios2_qsys_jtag_debug_module_write             (mm_interconnect_0_nios2_qsys_jtag_debug_module_write),       //                                         .write
		.nios2_qsys_jtag_debug_module_read              (mm_interconnect_0_nios2_qsys_jtag_debug_module_read),        //                                         .read
		.nios2_qsys_jtag_debug_module_readdata          (mm_interconnect_0_nios2_qsys_jtag_debug_module_readdata),    //                                         .readdata
		.nios2_qsys_jtag_debug_module_writedata         (mm_interconnect_0_nios2_qsys_jtag_debug_module_writedata),   //                                         .writedata
		.nios2_qsys_jtag_debug_module_byteenable        (mm_interconnect_0_nios2_qsys_jtag_debug_module_byteenable),  //                                         .byteenable
		.nios2_qsys_jtag_debug_module_waitrequest       (mm_interconnect_0_nios2_qsys_jtag_debug_module_waitrequest), //                                         .waitrequest
		.nios2_qsys_jtag_debug_module_debugaccess       (mm_interconnect_0_nios2_qsys_jtag_debug_module_debugaccess), //                                         .debugaccess
		.onchip_memory2_s1_address                      (mm_interconnect_0_onchip_memory2_s1_address),                //                        onchip_memory2_s1.address
		.onchip_memory2_s1_write                        (mm_interconnect_0_onchip_memory2_s1_write),                  //                                         .write
		.onchip_memory2_s1_readdata                     (mm_interconnect_0_onchip_memory2_s1_readdata),               //                                         .readdata
		.onchip_memory2_s1_writedata                    (mm_interconnect_0_onchip_memory2_s1_writedata),              //                                         .writedata
		.onchip_memory2_s1_byteenable                   (mm_interconnect_0_onchip_memory2_s1_byteenable),             //                                         .byteenable
		.onchip_memory2_s1_chipselect                   (mm_interconnect_0_onchip_memory2_s1_chipselect),             //                                         .chipselect
		.onchip_memory2_s1_clken                        (mm_interconnect_0_onchip_memory2_s1_clken),                  //                                         .clken
		.sysid_qsys_control_slave_address               (mm_interconnect_0_sysid_qsys_control_slave_address),         //                 sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata              (mm_interconnect_0_sysid_qsys_control_slave_readdata)         //                                         .readdata
	);

	esn7e_demo_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (nios2_qsys_d_irq_irq)            //    sender.irq
	);

	esn7e_demo_avalon_st_adapter #(
		.inBitsPerSymbol (32),
		.inUsePackets    (0),
		.inDataWidth     (32),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (0),
		.inReadyLatency  (0),
		.outDataWidth    (32),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (1)
	) avalon_st_adapter (
		.in_clk_0_clk   (altpll_esn_c0_clk),                                                // in_clk_0.clk
		.in_rst_0_reset (esn_reset_gate_reset_out_reset),                                   // in_rst_0.reset
		.in_0_valid     (echostatenetwork_7units_expanded_0_avalon_streaming_source_valid), //     in_0.valid
		.in_0_data      (echostatenetwork_7units_expanded_0_avalon_streaming_source_data),  //         .data
		.out_0_valid    (avalon_st_adapter_out_0_valid),                                    //    out_0.valid
		.out_0_data     (avalon_st_adapter_out_0_data),                                     //         .data
		.out_0_ready    (avalon_st_adapter_out_0_ready)                                     //         .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (nios2_qsys_jtag_debug_module_reset_reset), // reset_in0.reset
		.reset_in1      (~reset_reset_n),                           // reset_in1.reset
		.clk            (clk_clk),                                  //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),           // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),       //          .reset_req
		.reset_req_in0  (1'b0),                                     // (terminated)
		.reset_req_in1  (1'b0),                                     // (terminated)
		.reset_in2      (1'b0),                                     // (terminated)
		.reset_req_in2  (1'b0),                                     // (terminated)
		.reset_in3      (1'b0),                                     // (terminated)
		.reset_req_in3  (1'b0),                                     // (terminated)
		.reset_in4      (1'b0),                                     // (terminated)
		.reset_req_in4  (1'b0),                                     // (terminated)
		.reset_in5      (1'b0),                                     // (terminated)
		.reset_req_in5  (1'b0),                                     // (terminated)
		.reset_in6      (1'b0),                                     // (terminated)
		.reset_req_in6  (1'b0),                                     // (terminated)
		.reset_in7      (1'b0),                                     // (terminated)
		.reset_req_in7  (1'b0),                                     // (terminated)
		.reset_in8      (1'b0),                                     // (terminated)
		.reset_req_in8  (1'b0),                                     // (terminated)
		.reset_in9      (1'b0),                                     // (terminated)
		.reset_req_in9  (1'b0),                                     // (terminated)
		.reset_in10     (1'b0),                                     // (terminated)
		.reset_req_in10 (1'b0),                                     // (terminated)
		.reset_in11     (1'b0),                                     // (terminated)
		.reset_req_in11 (1'b0),                                     // (terminated)
		.reset_in12     (1'b0),                                     // (terminated)
		.reset_req_in12 (1'b0),                                     // (terminated)
		.reset_in13     (1'b0),                                     // (terminated)
		.reset_req_in13 (1'b0),                                     // (terminated)
		.reset_in14     (1'b0),                                     // (terminated)
		.reset_req_in14 (1'b0),                                     // (terminated)
		.reset_in15     (1'b0),                                     // (terminated)
		.reset_req_in15 (1'b0)                                      // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (nios2_qsys_jtag_debug_module_reset_reset), // reset_in0.reset
		.reset_in1      (~reset_reset_n),                           // reset_in1.reset
		.clk            (),                                         //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),       // reset_out.reset
		.reset_req      (),                                         // (terminated)
		.reset_req_in0  (1'b0),                                     // (terminated)
		.reset_req_in1  (1'b0),                                     // (terminated)
		.reset_in2      (1'b0),                                     // (terminated)
		.reset_req_in2  (1'b0),                                     // (terminated)
		.reset_in3      (1'b0),                                     // (terminated)
		.reset_req_in3  (1'b0),                                     // (terminated)
		.reset_in4      (1'b0),                                     // (terminated)
		.reset_req_in4  (1'b0),                                     // (terminated)
		.reset_in5      (1'b0),                                     // (terminated)
		.reset_req_in5  (1'b0),                                     // (terminated)
		.reset_in6      (1'b0),                                     // (terminated)
		.reset_req_in6  (1'b0),                                     // (terminated)
		.reset_in7      (1'b0),                                     // (terminated)
		.reset_req_in7  (1'b0),                                     // (terminated)
		.reset_in8      (1'b0),                                     // (terminated)
		.reset_req_in8  (1'b0),                                     // (terminated)
		.reset_in9      (1'b0),                                     // (terminated)
		.reset_req_in9  (1'b0),                                     // (terminated)
		.reset_in10     (1'b0),                                     // (terminated)
		.reset_req_in10 (1'b0),                                     // (terminated)
		.reset_in11     (1'b0),                                     // (terminated)
		.reset_req_in11 (1'b0),                                     // (terminated)
		.reset_in12     (1'b0),                                     // (terminated)
		.reset_req_in12 (1'b0),                                     // (terminated)
		.reset_in13     (1'b0),                                     // (terminated)
		.reset_req_in13 (1'b0),                                     // (terminated)
		.reset_in14     (1'b0),                                     // (terminated)
		.reset_req_in14 (1'b0),                                     // (terminated)
		.reset_in15     (1'b0),                                     // (terminated)
		.reset_req_in15 (1'b0)                                      // (terminated)
	);

endmodule
