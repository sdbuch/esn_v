module rdout_top(ce, sclr, sysclk, Q);

input ce, sclr, sysclk;
output [17:0] Q;


endmodule
