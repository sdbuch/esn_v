module pe_16x4_top(ce, sclr, sysclk, Q0, Q1, Q2, Q3);



endmodule
